module buffer(I, O);
	input I;
	output O;
	buf gate(O, I);
endmodule	