module half_adder(A,B,C,SUM);
input A,B;
output C, SUM;

xor x1(SUM, A,B);
and a1(C, A,B);
endmodule
